module SIPS4 (
	input wire clk // 50MHz input clock
);
endmodule